// niosII.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module niosII (
		input  wire  clk_clk,           //        clk.clk
		input  wire  reset_reset_n,     //      reset.reset_n
		input  wire  sem_export_train,  // sem_export.train
		output wire  sem_export_red,    //           .red
		output wire  sem_export_yellow, //           .yellow
		output wire  sem_export_green   //           .green
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [17:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [17:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sem_ctl_slave_readdata;                  // sem:ctl_rddata -> mm_interconnect_0:sem_ctl_slave_readdata
	wire   [1:0] mm_interconnect_0_sem_ctl_slave_address;                   // mm_interconnect_0:sem_ctl_slave_address -> sem:ctl_addr
	wire         mm_interconnect_0_sem_ctl_slave_read;                      // mm_interconnect_0:sem_ctl_slave_read -> sem:ctl_rd
	wire         mm_interconnect_0_sem_ctl_slave_write;                     // mm_interconnect_0:sem_ctl_slave_write -> sem:ctl_wr
	wire  [31:0] mm_interconnect_0_sem_ctl_slave_writedata;                 // mm_interconnect_0:sem_ctl_slave_writedata -> sem:ctl_wrdata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire   [1:0] mm_interconnect_0_sem_ram_slave_address;                   // mm_interconnect_0:sem_ram_slave_address -> sem:ram_addr
	wire         mm_interconnect_0_sem_ram_slave_write;                     // mm_interconnect_0:sem_ram_slave_write -> sem:ram_wr
	wire  [31:0] mm_interconnect_0_sem_ram_slave_writedata;                 // mm_interconnect_0:sem_ram_slave_writedata -> sem:ram_wrdata
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;             // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;               // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                  // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;              // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_mem_s2_chipselect;                       // mm_interconnect_0:mem_s2_chipselect -> mem:chipselect2
	wire  [31:0] mm_interconnect_0_mem_s2_readdata;                         // mem:readdata2 -> mm_interconnect_0:mem_s2_readdata
	wire  [14:0] mm_interconnect_0_mem_s2_address;                          // mm_interconnect_0:mem_s2_address -> mem:address2
	wire   [3:0] mm_interconnect_0_mem_s2_byteenable;                       // mm_interconnect_0:mem_s2_byteenable -> mem:byteenable2
	wire         mm_interconnect_0_mem_s2_write;                            // mm_interconnect_0:mem_s2_write -> mem:write2
	wire  [31:0] mm_interconnect_0_mem_s2_writedata;                        // mm_interconnect_0:mem_s2_writedata -> mem:writedata2
	wire         mm_interconnect_0_mem_s2_clken;                            // mm_interconnect_0:mem_s2_clken -> mem:clken2
	wire         mm_interconnect_0_mem_s1_chipselect;                       // mm_interconnect_0:mem_s1_chipselect -> mem:chipselect
	wire  [31:0] mm_interconnect_0_mem_s1_readdata;                         // mem:readdata -> mm_interconnect_0:mem_s1_readdata
	wire  [14:0] mm_interconnect_0_mem_s1_address;                          // mm_interconnect_0:mem_s1_address -> mem:address
	wire   [3:0] mm_interconnect_0_mem_s1_byteenable;                       // mm_interconnect_0:mem_s1_byteenable -> mem:byteenable
	wire         mm_interconnect_0_mem_s1_write;                            // mm_interconnect_0:mem_s1_write -> mem:write
	wire  [31:0] mm_interconnect_0_mem_s1_writedata;                        // mm_interconnect_0:mem_s1_writedata -> mem:writedata
	wire         mm_interconnect_0_mem_s1_clken;                            // mm_interconnect_0:mem_s1_clken -> mem:clken
	wire         irq_mapper_receiver0_irq;                                  // sys_clk_timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, mem:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sys_clk_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, mem:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [mm_interconnect_0:sem_reset_sink_reset_bridge_in_reset_reset, sem:clrn]

	niosII_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	niosII_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	niosII_mem mem (
		.address     (mm_interconnect_0_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_mem_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_mem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_mem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_mem_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_mem_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_mem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_mem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_mem_s2_byteenable), //       .byteenable
		.clk         (clk_clk),                             //   clk1.clk
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                 // (terminated)
	);

	dec #(
		.m (8)
	) sem (
		.clk        (clk_clk),                                   //      clock.clk
		.clrn       (~rst_controller_001_reset_out_reset),       // reset_sink.reset_n
		.ctl_wr     (mm_interconnect_0_sem_ctl_slave_write),     //  ctl_slave.write
		.ctl_rd     (mm_interconnect_0_sem_ctl_slave_read),      //           .read
		.ctl_addr   (mm_interconnect_0_sem_ctl_slave_address),   //           .address
		.ctl_wrdata (mm_interconnect_0_sem_ctl_slave_writedata), //           .writedata
		.ctl_rddata (mm_interconnect_0_sem_ctl_slave_readdata),  //           .readdata
		.ram_wr     (mm_interconnect_0_sem_ram_slave_write),     //  ram_slave.write
		.ram_addr   (mm_interconnect_0_sem_ram_slave_address),   //           .address
		.ram_wrdata (mm_interconnect_0_sem_ram_slave_writedata), //           .writedata
		.train      (sem_export_train),                          //        sem.train
		.red        (sem_export_red),                            //           .red
		.yellow     (sem_export_yellow),                         //           .yellow
		.green      (sem_export_green)                           //           .green
	);

	niosII_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                       //   irq.irq
	);

	niosII_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                (clk_clk),                                                   //                              clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                            //      cpu_reset_reset_bridge_in_reset.reset
		.sem_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // sem_reset_sink_reset_bridge_in_reset.reset
		.cpu_data_master_address                    (cpu_data_master_address),                                   //                      cpu_data_master.address
		.cpu_data_master_waitrequest                (cpu_data_master_waitrequest),                               //                                     .waitrequest
		.cpu_data_master_byteenable                 (cpu_data_master_byteenable),                                //                                     .byteenable
		.cpu_data_master_read                       (cpu_data_master_read),                                      //                                     .read
		.cpu_data_master_readdata                   (cpu_data_master_readdata),                                  //                                     .readdata
		.cpu_data_master_write                      (cpu_data_master_write),                                     //                                     .write
		.cpu_data_master_writedata                  (cpu_data_master_writedata),                                 //                                     .writedata
		.cpu_data_master_debugaccess                (cpu_data_master_debugaccess),                               //                                     .debugaccess
		.cpu_instruction_master_address             (cpu_instruction_master_address),                            //               cpu_instruction_master.address
		.cpu_instruction_master_waitrequest         (cpu_instruction_master_waitrequest),                        //                                     .waitrequest
		.cpu_instruction_master_read                (cpu_instruction_master_read),                               //                                     .read
		.cpu_instruction_master_readdata            (cpu_instruction_master_readdata),                           //                                     .readdata
		.cpu_debug_mem_slave_address                (mm_interconnect_0_cpu_debug_mem_slave_address),             //                  cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                  (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                     .write
		.cpu_debug_mem_slave_read                   (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                     .read
		.cpu_debug_mem_slave_readdata               (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                     .readdata
		.cpu_debug_mem_slave_writedata              (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                     .writedata
		.cpu_debug_mem_slave_byteenable             (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                     .byteenable
		.cpu_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                     .waitrequest
		.cpu_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                     .debugaccess
		.jtag_uart_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                     .write
		.jtag_uart_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                     .read
		.jtag_uart_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                     .chipselect
		.mem_s1_address                             (mm_interconnect_0_mem_s1_address),                          //                               mem_s1.address
		.mem_s1_write                               (mm_interconnect_0_mem_s1_write),                            //                                     .write
		.mem_s1_readdata                            (mm_interconnect_0_mem_s1_readdata),                         //                                     .readdata
		.mem_s1_writedata                           (mm_interconnect_0_mem_s1_writedata),                        //                                     .writedata
		.mem_s1_byteenable                          (mm_interconnect_0_mem_s1_byteenable),                       //                                     .byteenable
		.mem_s1_chipselect                          (mm_interconnect_0_mem_s1_chipselect),                       //                                     .chipselect
		.mem_s1_clken                               (mm_interconnect_0_mem_s1_clken),                            //                                     .clken
		.mem_s2_address                             (mm_interconnect_0_mem_s2_address),                          //                               mem_s2.address
		.mem_s2_write                               (mm_interconnect_0_mem_s2_write),                            //                                     .write
		.mem_s2_readdata                            (mm_interconnect_0_mem_s2_readdata),                         //                                     .readdata
		.mem_s2_writedata                           (mm_interconnect_0_mem_s2_writedata),                        //                                     .writedata
		.mem_s2_byteenable                          (mm_interconnect_0_mem_s2_byteenable),                       //                                     .byteenable
		.mem_s2_chipselect                          (mm_interconnect_0_mem_s2_chipselect),                       //                                     .chipselect
		.mem_s2_clken                               (mm_interconnect_0_mem_s2_clken),                            //                                     .clken
		.sem_ctl_slave_address                      (mm_interconnect_0_sem_ctl_slave_address),                   //                        sem_ctl_slave.address
		.sem_ctl_slave_write                        (mm_interconnect_0_sem_ctl_slave_write),                     //                                     .write
		.sem_ctl_slave_read                         (mm_interconnect_0_sem_ctl_slave_read),                      //                                     .read
		.sem_ctl_slave_readdata                     (mm_interconnect_0_sem_ctl_slave_readdata),                  //                                     .readdata
		.sem_ctl_slave_writedata                    (mm_interconnect_0_sem_ctl_slave_writedata),                 //                                     .writedata
		.sem_ram_slave_address                      (mm_interconnect_0_sem_ram_slave_address),                   //                        sem_ram_slave.address
		.sem_ram_slave_write                        (mm_interconnect_0_sem_ram_slave_write),                     //                                     .write
		.sem_ram_slave_writedata                    (mm_interconnect_0_sem_ram_slave_writedata),                 //                                     .writedata
		.sys_clk_timer_s1_address                   (mm_interconnect_0_sys_clk_timer_s1_address),                //                     sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                     (mm_interconnect_0_sys_clk_timer_s1_write),                  //                                     .write
		.sys_clk_timer_s1_readdata                  (mm_interconnect_0_sys_clk_timer_s1_readdata),               //                                     .readdata
		.sys_clk_timer_s1_writedata                 (mm_interconnect_0_sys_clk_timer_s1_writedata),              //                                     .writedata
		.sys_clk_timer_s1_chipselect                (mm_interconnect_0_sys_clk_timer_s1_chipselect)              //                                     .chipselect
	);

	niosII_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
